module HA (
  input A, B,
  output S, C
);


endmodule